edit on web
