package test_pkg;

  import counter_pkg::*;

  `include "base_test.sv"
  `include "count_up_test.sv"
  `include "count_down_test.sv"
  `include "count_down_with_data_test.sv"
  `include "count_up_with_data_test.sv"
endpackage
