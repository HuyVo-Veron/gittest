package src_snk_pkg;

  `include "packet.sv"
  `include "source.sv"
  `include "sink.sv"

endpackage
