class packet;
	int pid;

	function new(int i);
		pid = i;
	endfunction

endclass

