package apb_pkg;
  import uvm_pkg::*;

  `include "apb_transaction.sv"
  `include "apb_sequencer.sv"
  `include "apb_driver.sv"
  `include "apb_monitor.sv"
  `include "apb_agent.sv"
endpackage: apb_pkg
