import uvm_pkg::*;
import ahb_pkg::*;

module testbench;

  initial begin
    /** Start the UVM test */
    run_test();
  end

endmodule

