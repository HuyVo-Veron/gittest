package counter_pkg;

  `include "packet.sv"
  `include "stimulus.sv"
  `include "driver.svp"
  `include "monitor.svp"
  `include "scoreboard.sv"
  `include "environment.sv"

endpackage
