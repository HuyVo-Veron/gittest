import uvm_pkg::*;
import apb_pkg::*;

module testbench;

  initial begin
    /** Start the UVM test */
    run_test();
  end

endmodule

