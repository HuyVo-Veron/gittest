interface dut_if;
  logic       clk;
  logic       rst_n;
  logic       valid;
  logic[7:0]  data_in;
  logic       TXD;

endinterface
