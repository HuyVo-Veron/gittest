package ahb_pkg;
  import uvm_pkg::*;

  `include "ahb_transaction.sv"
  `include "ahb_sequencer.sv"
  `include "ahb_driver.sv"
  `include "ahb_monitor.sv"
  `include "ahb_agent.sv"
endpackage: ahb_pkg
