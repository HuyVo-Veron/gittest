edit on web

add from vnc

