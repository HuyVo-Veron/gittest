package data_type_pkg;
	typedef struct{
		bit [2:0] pid;
		bit [7:0] data;
		} packet_st;

endpackage
